module top_module(
    input [31:0] a,
    input [31:0] b,
    
    output [31:0] sum
);
    wire cin, cout1, cout2;
    assign cin = 0;
    add16 inst1(.a(a[15:0]), .b(b[15:0]), .cin(cin), .sum(sum[15:0]), .cout(cout1));
    add16 inst2(.a(a[31:16]), .b(b[31:16]), .cin(cout1), .sum(sum[31:16]), .cout(cout2));
endmodule
